module wallace(a,b,c0,c1);

	input [52:0] a,b;
	wire [0:211] c;
	
	output [0:105] c0,c1;
	
	wire [0:5617] u;
	wire [0:2861] u1;
	wire [0:1271] u2;
	wire [0:635] u3;
	wire [0:635] u4;
	wire [0:317] u5; 
	
	partialProductGenerator pp(a,b,u);
	
	
	c16 #(0) c161(u[0:635],u1[0:317]);
	c16 #(6) c162(u[636:1271],u1[318:635]);
	c16 #(12) c163(u[1272:1907],u1[636:953]);
	c16 #(18) c164(u[1906:2543],u1[954:1271]);
	c16 #(24) c165(u[2542:3179],u1[1272:1589]);
	c16 #(30) c166(u[3180:3815],u1[1590:1907]);
	c16 #(36) c167(u[3816:4451],u1[1908:2225]);
	c16 #(42) c168(u[4452:5087],u1[2226:2543]);
	c5 #(0) c51(u[5088:5617],u1[2544:2861]);
	
	c26 #(0) c261(u1[0:635],u2[0:317]);
	c26 #(12) c262(u1[636:1271],u2[318:635]);
	c26 #(24) c263(u1[1272:1907],u2[636:953]);
	c26 #(36) c264(u1[1906:2543],u2[954:1271]);
	
	c36 #(0) c361(u2[0:635],u3[0:317]);
	c36 #(24) c362(u2[636:1271],u3[318:635]);
	
	c46 #(0) c461(u3[0:635],u4[0:317]);
	
	assign u4[318:635]=u1[2544:2861];
	
	c56 #(0) c561(u4[0:635],u5[0:317]);
	
	c3 #(0) c31 (u5[0:317],c[0:211]);
	
	assign c0[0:105]=c[0:105];
	assign c1[0:105]=c[106:211];
	/*
	always@(posedge clk)
	begin
		ur<=u;
	end
	
	initial
	begin
		assign u=5618'b0;
		assign u1=2862'b0;
		assign u2=1272'b0;
		assign u3=636'b0;
		assign u4=636'b0;
		assign u5=318'b0;
		assign c=212'b0;	
	end
*/
endmodule
